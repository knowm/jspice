* Qucs 0.0.19  /Users/marendall/.qucs/KnowmMemristor_prj/knowm_mr_pulse.sch
VPr1 Vin Vmr DC 0
R1 0 Vout  500

YMEMRISTOR MR1 Vmr  Vout MRM5
V1 Vin 0 DC 0 PULSE( 2  0 0N 1N 1N 5e-06 1.0002e-05)  AC 0
.model MRM5 memristor ( level=5
+ Roff=1500 Ron=500 Voff=0.27 Von=0.27
+ Tau=0.0001 Phi=1.0
+ Sfa=0.0 Sfb=0.0 Sra=0.0 Srb=0.0  Rinit=500 )

.STEP V1:V2 LIST 0.25 0.5 0.75 1.0
.tran 1us 50us
.PRINT  tran format=raw file=knowm_mr_pulse_tran.txt I(VPr1) v(Vin) v(Vmr) v(Vout)
.END
